library verilog;
use verilog.vl_types.all;
entity switch_vlg_tst is
end switch_vlg_tst;
